-------------------------------------------------------------------------------
--
-- Title       : No Title
-- Design      : top_level
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : U:\workspace\nexysterm\Aldec\compile\vga_top.vhd
-- Generated   : Wed Jul  4 18:26:49 2012
-- From        : U:\workspace\nexysterm\Aldec\src\vga_top.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library unisim;
use unisim.vcomponents.all;
use work.VGA_TIMING.all;

entity vga_top is
    port(
        i_sys_reset : in STD_LOGIC;
        i_tram_clk : in STD_LOGIC;
        i_tram_en : in STD_LOGIC;
        i_tram_addr : in STD_LOGIC_VECTOR(10 downto 0);
        i_tram_data : in STD_LOGIC_VECTOR(15 downto 0);
        i_vga_clk : in STD_LOGIC;
        o_vga_hsync : out STD_LOGIC;
        o_vga_vsync : out STD_LOGIC;
        o_vga_blu : out STD_LOGIC_VECTOR(1 downto 0);
        o_vga_grn : out STD_LOGIC_VECTOR(2 downto 0);
        o_vga_red : out STD_LOGIC_VECTOR(2 downto 0)
    );
end vga_top;

architecture vga_top of vga_top is
---- Component declarations -----
component char_rom
    port (
        CLK : in STD_LOGIC;
        i_char : in STD_LOGIC_VECTOR(7 downto 0);
        i_col : in STD_LOGIC_VECTOR(2 downto 0);
        i_row : in STD_LOGIC_VECTOR(3 downto 0);
        o_bit : out STD_LOGIC
    );
end component;
component text_ram
    port (
        i_rd_addr : in STD_LOGIC_VECTOR(10 downto 0);
        i_rd_clk : in STD_LOGIC;
        i_wr_addr : in STD_LOGIC_VECTOR(10 downto 0);
        i_wr_clk : in STD_LOGIC;
        i_wr_data : in STD_LOGIC_VECTOR(15 downto 0);
        i_wr_en : in STD_LOGIC;
        o_rd_data : out STD_LOGIC_VECTOR(15 downto 0)
    );
end component;
component VGA_Timer
    port (
        ref_clk : in STD_LOGIC;
        reset : in STD_LOGIC;
        o_chrx : out INTEGER range 79 downto 0;
        o_chry : out INTEGER range 39 downto 0;
        o_schrx : out INTEGER range 7 downto 0;
        o_schry : out INTEGER range 11 downto 0;
        o_x_blank : out STD_LOGIC;
        o_x_pos : out INTEGER range H_TOTAL-1 downto 0;
        o_x_sync : out STD_LOGIC;
        o_y_blank : out STD_LOGIC;
        o_y_pos : out INTEGER range V_TOTAL-1 downto 0;
        o_y_sync : out STD_LOGIC
    );
end component;

---- Signal declarations used on the diagram ----
--signal s_bit : STD_LOGIC;
--signal s_chrx : INTEGER range 79 downto 0;
--signal s_chry : INTEGER range 39 downto 0;
--signal s_hsync : STD_LOGIC;
--signal s_schrx : INTEGER range 7 downto 0;
--signal s_schry : INTEGER range 11 downto 0;
--signal s_vsync : STD_LOGIC;
--signal s_xblank : STD_LOGIC;
--signal s_xpos : INTEGER range H_TOTAL-1 downto 0;
--signal s_xsync : STD_LOGIC;
--signal s_yblank : STD_LOGIC;
--signal s_ypos : INTEGER range V_TOTAL-1 downto 0;
--signal s_ysync : STD_LOGIC;
--signal s_blu : STD_LOGIC_VECTOR (1 downto 0);
--signal s_char : STD_LOGIC_VECTOR (15 downto 0);
--signal s_col : STD_LOGIC_VECTOR (2 downto 0);
--signal s_grn : STD_LOGIC_VECTOR (2 downto 0);
--signal s_rd_addr : STD_LOGIC_VECTOR (10 downto 0);
--signal s_red : STD_LOGIC_VECTOR (2 downto 0);
--signal s_row : STD_LOGIC_VECTOR (3 downto 0);

-- VGA Timer output signals
signal s_tmr_chrx    : integer range 79 downto 0;
signal s_tmr_chry    : integer range 39 downto 0;
signal s_tmr_schrx   : integer range 7 downto 0;
signal s_tmr_schry   : integer range 11 downto 0;
signal s_tmr_x_blank : std_logic;
signal s_tmr_y_blank : std_logic;
signal s_tmr_x_sync  : std_logic;
signal s_tmr_y_sync  : std_logic;

signal s_rd_addr : std_logic_vector(10 downto 0);

-- TRAM output signals
signal s_tram_x_blank : std_logic;
signal s_tram_y_blank : std_logic;
signal s_tram_x_sync  : std_logic;
signal s_tram_y_sync  : std_logic;
signal s_tram_row   : std_logic_vector(3 downto 0);
signal s_tram_col   : std_logic_vector(2 downto 0);
signal s_tram_data  : std_logic_vector(15 downto 0);
signal s_tram_char  : std_logic_vector(7 downto 0);

-- CROM output signals
signal s_crom_x_blank : std_logic;
signal s_crom_y_blank : std_logic;
signal s_crom_x_sync  : std_logic;
signal s_crom_y_sync  : std_logic;
signal s_crom_color   : std_logic_vector(7 downto 0);
signal s_crom_bit     : std_logic;


begin

vga_timer_inst : VGA_Timer
    port map(
        ref_clk     => i_vga_clk,
        reset       => i_sys_reset,
        
        o_x_pos     => open,
        o_y_pos     => open,
        
        o_chrx      => s_tmr_chrx,
        o_chry      => s_tmr_chry,
        
        o_schrx     => s_tmr_schrx,
        o_schry     => s_tmr_schry,
        
        o_x_blank   => s_tmr_x_blank,
        o_y_blank   => s_tmr_y_blank,
        o_x_sync    => s_tmr_x_sync,
        o_y_sync    => s_tmr_y_sync
    );

-- ----------

s_rd_addr <= std_logic_vector(to_unsigned((s_tmr_chrx + (100*s_tmr_chry)),s_rd_addr'length));

tram_inst : text_ram
    port map(
        i_rd_clk => i_vga_clk,
        i_rd_addr => s_rd_addr,
        o_rd_data => s_tram_data,
        
        i_wr_addr => i_tram_addr,
        i_wr_clk => i_tram_clk,
        i_wr_data => i_tram_data,
        i_wr_en => i_tram_en
    );

-- Delay everything that didn't go through the TRAM
process(i_vga_clk) begin
    if rising_edge(i_vga_clk) then
        s_tram_col <= std_logic_vector(to_unsigned(s_tmr_schrx,s_tram_col'length));
        s_tram_row <= std_logic_vector(to_unsigned(s_tmr_schry,s_tram_row'length));
        s_tram_x_blank <= s_tmr_x_blank;
        s_tram_y_blank <= s_tmr_y_blank;
        s_tram_x_sync  <= s_tmr_x_sync;
        s_tram_y_sync  <= s_tmr_y_sync;
    end if;
end process;

-- ----------

s_tram_char <= s_tram_data(7 downto 0);

crom_inst : char_rom
    port map(
        CLK => i_vga_clk,
        i_char => s_tram_char,
        i_col => s_tram_col,
        i_row => s_tram_row,
        o_bit => s_crom_bit
    );

-- Delay everything that didn't go through the CROM
process(i_vga_clk) begin
    if rising_edge(i_vga_clk) then
        s_crom_color <= s_tram_data(15 downto 8);
        s_crom_x_blank <= s_tram_x_blank;
        s_crom_y_blank <= s_tram_y_blank;
        s_crom_x_sync  <= s_tram_x_sync;
        s_crom_y_sync  <= s_tram_y_sync;
    end if;
end process;

-- ----------

process (i_vga_clk) begin
    if rising_edge(i_vga_clk) then
        o_vga_hsync <= s_crom_x_sync;
        o_vga_vsync <= s_crom_y_sync;
        if (s_crom_x_blank='0' and s_crom_y_blank='0' and s_crom_bit='1') then
            o_vga_red <= s_crom_color(7 downto 5);
            o_vga_grn <= s_crom_color(4 downto 2);
            o_vga_blu <= s_crom_color(1 downto 0);
        else
            o_vga_red <= (others => '0');
            o_vga_grn <= (others => '0');
            o_vga_blu <= (others => '0');
        end if;
    end if;
end process;

end vga_top;
