----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:06:45 07/01/2012 
-- Design Name: 
-- Module Name:    CRG - behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
use UNISIM.VComponents.all;

entity char_rom is
    Port (
        CLK : in  std_logic;
        --i_reset : in  std_logic;
        
        i_char : in std_logic_vector(7 downto 0);
        i_col : in std_logic_vector(2 downto 0);
        i_row : in std_logic_vector(3 downto 0);
        
        o_bit : out std_logic
    );
end char_rom;

architecture Behavioral of char_rom is
    signal DO1, DO2 : std_logic_vector(0 downto 0);
    signal FULL_ADDR : std_logic_vector(14 downto 0);
    signal ADDR : std_logic_vector(13 downto 0);
begin
    FULL_ADDR <= i_char & i_row & i_col;
    ADDR <= FULL_ADDR(13 downto 0);
    
    o_bit <= DO1(0) when FULL_ADDR(14)='0' else DO2(0);

char_rom_bram1 : RAMB16_S1
    generic map (
        INIT => X"0", -- Value of output RAM registers at startup
        SRVAL => X"0", -- Ouput value upon SSR assertion
        WRITE_MODE => "WRITE_FIRST", -- WRITE_FIRST, READ_FIRST or NO_CHANGE
INIT_00 => X"00000000000000003b6e003b6e00000000000000007ee7e7ffe7e7cf9999c37e",
INIT_01 => X"00000000000076db1bfbdbdb76000000000000000000761b1b1b7b1b1b1b1b76",
INIT_02 => X"0000000000101010107c0011111f111100000000000000081c3e7f3e1c080000",
INIT_03 => X"000000000044247c443c001e0101011e000000000004041c047c00010107011f",
INIT_04 => X"00000000114411441144114411441144000000000004041c047c001f01010101",
INIT_05 => X"00000000dd77dd77dd77dd77dd77dd770000000055aa55aa55aa55aa55aa55aa",
INIT_06 => X"00000000ffffffffffff00000000000000000000ffffffffffffffffffffffff",
INIT_07 => X"000000000f0f0f0f0f0f0f0f0f0f0f0f00000000000000000000ffffffffffff",
INIT_08 => X"00000000007c0404040400111915131100000000f0f0f0f0f0f0f0f0f0f0f0f0",
INIT_09 => X"000000000000007e007e0c18306000000000000000101010107c00040a0a1111",
INIT_0a => X"0000000000000003067f1c7f30600000000000000000007e007e30180c060000",
INIT_0b => X"00000000000001070f3f7f3f0f07010000000000000040707c7e7f7e7c704000",
INIT_0c => X"000000000000183c7e181818181818000000000000001818181818187e3c1800",
INIT_0d => X"00000000000000000c067f060c000000000000000000000018307f3018000000",
INIT_0e => X"000000000000000014367f3614000000000000000000183c7e1818187e3c1800",
INIT_0f => X"00000000000000363636763e0300000000000000000000000c067f666c606000",
INIT_10 => X"00000000000018180018183c3c3c180000000000000000000000000000000000",
INIT_11 => X"000000000000367f3636367f36000000000000000000000000000000286c6c00",
INIT_12 => X"00000000000063660c18306646000000000000000000083e6b381c0e6b3e0800",
INIT_13 => X"000000000000000000000000183038380000000000006e33337f4e1c1c361c00",
INIT_14 => X"0000000000000c183030303030180c0000000000000030180c0c0c0c0c183000",
INIT_15 => X"000000000000000018187e18180000000000000000000000361c7f1c36000000",
INIT_16 => X"000000000000000000007f000000000000000000001830303000000000000000",
INIT_17 => X"0000000000000003060c18306000000000000000000018180000000000000000",
INIT_18 => X"0000000000007e1818181818181e18000000000000003e6363636b6363633e00",
INIT_19 => X"0000000000003e6360603c6060633e000000000000007f63060c183063633e00",
INIT_1a => X"0000000000003e6360603f0303037f000000000000003030307f33363c383000",
INIT_1b => X"0000000000000c0c0c0c0c1830637f000000000000003e6363633f0303633e00",
INIT_1c => X"0000000000003e6360607e6363633e000000000000003e6363633e6363633e00",
INIT_1d => X"0000000000183030300000303000000000000000000000303000003030000000",
INIT_1e => X"0000000000000000007f007f0000000000000000000030180c0603060c183000",
INIT_1f => X"00000000000018180018183063633e00000000000000060c18306030180c0600",
INIT_20 => X"0000000000006363637f636363361c000000000000007e033b7b7b7b63633e00",
INIT_21 => X"0000000000003c660303030303663c000000000000003f6666663e6666663f00",
INIT_22 => X"0000000000007f6606063e0606667f000000000000001f366666666666361f00",
INIT_23 => X"0000000000003e636373030363633e000000000000000f0606063e0606667f00",
INIT_24 => X"0000000000003c181818181818183c00000000000000636363637f6363636300",
INIT_25 => X"0000000000006363331b0f0f1b3363000000000000000e1b1b18181818183c00",
INIT_26 => X"00000000000063636b6b6b7f776363000000000000007f664606060606060f00",
INIT_27 => X"0000000000003e636363636363633e000000000000006373737b6f6767636300",
INIT_28 => X"0000000000603e6b6363636363633e000000000000000f0606063e6666663f00",
INIT_29 => X"0000000000003e6360301c0603633e000000000000006766361e3e6666663f00",
INIT_2a => X"0000000000003e6363636363636363000000000000003c1818181818185a7e00",
INIT_2b => X"0000000000006363777f6b6b6b636300000000000000081c3663636363636300",
INIT_2c => X"0000000000003c1818183c66666666000000000000006363361c1c1c36636300",
INIT_2d => X"0000000000003e060606060606063e000000000000007f6343060c1831637f00",
INIT_2e => X"0000000000003e303030303030303e00000000000000006030180c0603000000",
INIT_2f => X"00000000ff0000000000000000000000000000000000000000000000663c1800",
INIT_30 => X"0000000000006e3b333e301e0000000000000000000000000000000030183838",
INIT_31 => X"0000000000003e630303633e000000000000000000003f666666663e06060700",
INIT_32 => X"0000000000003e63037f633e000000000000000000007e333333333e30303800",
INIT_33 => X"000000003e63607e6363736e000000000000000000001e0c0c0c3f0c0c6c3800",
INIT_34 => X"0000000000003c181818181c00181800000000000000676666666e3606060700",
INIT_35 => X"0000000000006766361e366606060700000000001e3333303030380030300000",
INIT_36 => X"00000000000063636b6b7f3600000000000000000000182c0c0c0c0c0c0c0e00",
INIT_37 => X"0000000000003e636363633e0000000000000000000066666666663b00000000",
INIT_38 => X"000000007830303e3333336e00000000000000000f06063e6666663b00000000",
INIT_39 => X"0000000000003e63380e633e000000000000000000000f060606663b00000000",
INIT_3a => X"0000000000006e333333333300000000000000000000386c0c0c0c3f0c0c0c00",
INIT_3b => X"000000000000367f6b6b636300000000000000000000081c3663636300000000",
INIT_3c => X"000000003e63606e736363630000000000000000000063361c1c366300000000",
INIT_3d => X"000000000000701818180e18181870000000000000007f460c18317f00000000",
INIT_3e => X"0000000000000e181818701818180e0000000000000018181818181818181800",
INIT_3f => X"0000000000003c18183c666666006666000000000000000000000000003b6e00"
    )
    port map (
        DO   => DO1,   -- 1-bit Data Output
        ADDR => ADDR, -- 14-bit Address Input
        CLK  => CLK,  -- Clock
        DI   => (others => '0'),   -- 1-bit Data Input
        EN   => '1',   -- RAM Enable Input
        SSR  => '0',  -- Synchronous Set/Reset Input
        WE   => '0'   -- Write Enable Input
    );

char_rom_bram2 : RAMB16_S1
    generic map (
        INIT => X"0", -- Value of output RAM registers at startup
        SRVAL => X"0", -- Ouput value upon SSR assertion
        WRITE_MODE => "WRITE_FIRST", -- WRITE_FIRST, READ_FIRST or NO_CHANGE
INIT_00 => X"00000000000063637f6363361c000c1800000000000063637f6363361c00180c",
INIT_01 => X"00000000000063637f6363361c003b6e00000000000063637f63633e001c361c",
INIT_02 => X"00000000000063637f63633e001c361c00000000000063637f6363361c003636",
INIT_03 => X"000000001c33183c6663030303663c000000000000007b1b1b1b7f1b1b1b1b7e",
INIT_04 => X"0000000000007f66063e06667f000c180000000000007f66063e06667f003018",
INIT_05 => X"0000000000007f66063e06667f0036360000000000007f66063e06667f00361c",
INIT_06 => X"0000000000003c18181818183c000c180000000000003c18181818183c003018",
INIT_07 => X"0000000000003c18181818183c0066660000000000003c18181818183c00663c",
INIT_08 => X"0000000000006363737b6f6763003b6e0000000000001f3666666f6666361f00",
INIT_09 => X"0000000000003e63636363633e000c180000000000003e63636363633e00180c",
INIT_0a => X"0000000000003e63636363633e003b6e0000000000003e63636363633e00361c",
INIT_0b => X"0000000000000000361c1c36000000000000000000003e63636363633e003636",
INIT_0c => X"0000000000003e63636363636300180c0000000000003f63676f6b7b73637e00",
INIT_0d => X"0000000000003e63636363636300361c0000000000003e636363636363000c18",
INIT_0e => X"0000000000003c18183c6666660018300000000000003e636363636363003636",
INIT_0f => X"0000000000013b6b6363336363633e000000000000000f063e6666663e060f00",
INIT_10 => X"00000000183c3c3c181800181800000000000000007f41000000000000000000",
INIT_11 => X"000000000000366f66060f0606361c00000000000000083e6b0b0b6b3e080000",
INIT_12 => X"00000000000018183c187e183c6666000000000000003c46061f061f06463c00",
INIT_13 => X"000000003e6363303e63633e0663633e0000000000003e63603e03633e001c36",
INIT_14 => X"0000000000007e8199a58585a599817e0000000000003e63380e633e001c3600",
INIT_15 => X"00000000000000006c361b366c000000000000000000000000007e007c36363c",
INIT_16 => X"000000000000000000007e0000000000000000000000006060607e0000000000",
INIT_17 => X"000000000000000000000000000000ff0000000000007e81a5a59da5a59d817e",
INIT_18 => X"0000000000007e0018187e18180000000000000000000000000000001c361c00",
INIT_19 => X"000000000000000000001c3618361c00000000000000000000003e0c18361c00",
INIT_1a => X"0000000003036f3333333333000000000000000000007f63461c30637f001c36",
INIT_1b => X"00000000000000000018180000000000000000000000d8d8d8d8dedbdbdbfe00",
INIT_1c => X"000000000000000000001e0c0c0e0c000000000000007f460c18317f001c3600",
INIT_1d => X"00000000000000001b366c361b000000000000000000000000003e001c36361c",
INIT_1e => X"000000000000365b1b7b5b360000000000000000000076fb9b1b1bfbdbdb7600",
INIT_1f => X"000000003e6363060c0c000c0c0000000000000000003c1818183c6666006666",
INIT_20 => X"0000000000000000000018181818181800000000000000000000000000ff0000",
INIT_21 => X"00000000000000000000f8181818181800000000000000000000f80000000000",
INIT_22 => X"0000000018181818181818181818181800000000181818181818180000000000",
INIT_23 => X"00000000181818181818f8181818181800000000181818181818f80000000000",
INIT_24 => X"000000000000000000001f1818181818000000000000000000001f0000000000",
INIT_25 => X"00000000000000000000ff181818181800000000000000000000ff0000000000",
INIT_26 => X"000000001818181818181f1818181818000000001818181818181f0000000000",
INIT_27 => X"00000000181818181818ff181818181800000000181818181818ff0000000000",
INIT_28 => X"0000000000000000003e3636363636360000000000000000ff00000000000000",
INIT_29 => X"000000000000000000fe06f636363636000000000000000000fc0cfc00000000",
INIT_2a => X"0000000036363636363636363636363600000000363636363636363e00000000",
INIT_2b => X"000000003636363636f606f636363636000000003636363636f606fe00000000",
INIT_2c => X"0000000000000000003f3037363636360000000000000000003f303f00000000",
INIT_2d => X"000000000000000000ff00f736363636000000000000000000ff00ff00000000",
INIT_2e => X"0000000036363636363730373636363600000000363636363637303f00000000",
INIT_2f => X"000000003636363636f700f736363636000000003636363636f700ff00000000",
INIT_30 => X"0000000000006e3b333e301e00060c180000000000006e3b333e301e00180c06",
INIT_31 => X"0000000000006e3b333e301e003b6e000000000000006e3b333e301e00331e0c",
INIT_32 => X"0000000000006e3b333e301e001c361c0000000000006e3b333e301e00363600",
INIT_33 => X"000000001c36183e630303633e0000000000000000007edb1bfed8db7e000000",
INIT_34 => X"0000000000003e63037f633e000c18300000000000003e63037f633e0030180c",
INIT_35 => X"0000000000003e63037f633e003636000000000000003e63037f633e00361c08",
INIT_36 => X"0000000000003c181818181c000c18300000000000003c181818181c00180c06",
INIT_37 => X"0000000000003c181818181c003636000000000000003c181818181c00663c18",
INIT_38 => X"00000000000066666666663b003b6e000000000000003e636363637e301e0c1e",
INIT_39 => X"0000000000003e636363633e000c18300000000000003e636363633e00180c06",
INIT_3a => X"0000000000003e636363633e003b6e000000000000003e636363633e00361c08",
INIT_3b => X"000000000000001818007e00181800000000000000003e636363633e00363600",
INIT_3c => X"0000000000006e3333333333000c06030000000000003f676f7b737e00000000",
INIT_3d => X"0000000000006e333333333300331e0c0000000000006e3333333333000c1830",
INIT_3e => X"000000003e63606e73636363000c18300000000000006e333333333300333300",
INIT_3f => X"000000003e63606e7363636300636300000000000f06061e3636361e06060f00"
    )
    port map (
        DO   => DO2,   -- 1-bit Data Output
        ADDR => ADDR, -- 14-bit Address Input
        CLK  => CLK,  -- Clock
        DI   => (others => '0'),   -- 1-bit Data Input
        EN   => '1',   -- RAM Enable Input
        SSR  => '0',  -- Synchronous Set/Reset Input
        WE   => '0'   -- Write Enable Input
    );


end architecture;
